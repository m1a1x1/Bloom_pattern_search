// Filenames for simulating:
//
`define DATA_FNAME      "example_data"
`define SETTINGS_FNAME  "example_settings"
`define OUTDATA_FNAME   "out_data"

// Bloom-filter parameters
//
`define MIN_S       4
`define MAX_S       16
`define HASH_CNT    10
`define HASH_WIDTH  12
